// This file is public domain, it can be freely copied without restrictions.
// SPDX-License-Identifier: CC0-1.0
// Adder DUT
`timescale 1ns/1ps

module packed_unpacked (
  input  [4:0] vec_i,
  input  [4:0][3:0] matrix_i,
  input  unpack_i [4:0],
  input  [3:0] vec_unpack_i [4:0],
  output out_o
);


endmodule
